module Top_Level(

input wire a,
output wire b

);

assign a = b;
endmodule

module b
(
	input wire clk,
	input wire n_rst
);
endmodule
